
module mux3to1(a,sel,out);

input a[3:0];  // declaring inputs for mux
input sel[1:0];  //declaring inputs for select 
output out;  // declaring output  


reg       out; // declaring into reg
wire[1:0] sel;
wire[3:0] a; // declaring wires to be used


always @( sel or a )  //initialising  always 
begin
   if( sel == 2'b00) 
      out = a[0]; 

   if( sel == 2'b01) 
      out = a[1];

   if( sel == 2'b10) 
      out = a[2];

   if( sel == 2'b11) 
      out = 1'bx;
end 

endmodule